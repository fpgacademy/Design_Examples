

module DE10_Standard_NiosVg_Computer
//=======================================================
//  PARAMETER declarations
//=======================================================
// #(
// )


//=======================================================
//  PORT declarations
//=======================================================
(
////////////////////////////////////
// FPGA Pins
////////////////////////////////////

// Clock pins
input               CLOCK_50,
input               CLOCK2_50,
input               CLOCK3_50,
input               CLOCK4_50,

// ADC
output              ADC_CONVST,
output              ADC_SCLK,
output              ADC_SDI,
input               ADC_SDO,

// Audio
input               AUD_ADCDAT,
inout               AUD_ADCLRCK,
inout               AUD_BCLK,
output              AUD_DACDAT,
inout               AUD_DACLRCK,
output              AUD_XCK,

// SDRAM
output      [12: 0] DRAM_ADDR,
output      [ 1: 0] DRAM_BA,
output              DRAM_CAS_N,
output              DRAM_CKE,
output              DRAM_CLK,
output              DRAM_CS_N,
inout       [15: 0] DRAM_DQ,
output              DRAM_LDQM,
output              DRAM_RAS_N,
output              DRAM_UDQM,
output              DRAM_WE_N,

// I2C Bus for Configuration of the Audio and Video-In Chips
output              FPGA_I2C_SCLK,
inout               FPGA_I2C_SDAT,

// 40-pin headers
inout       [35: 0] GPIO,

// Seven Segment Displays
output      [ 6: 0] HEX0,
output      [ 6: 0] HEX1,
output      [ 6: 0] HEX2,
output      [ 6: 0] HEX3,
output      [ 6: 0] HEX4,
output      [ 6: 0] HEX5,

// IR
input               IRDA_RXD,
output              IRDA_TXD,

// Pushbuttons
input       [ 3: 0] KEY,

// LEDs
output      [ 9: 0] LEDR,

// PS2 Ports
inout               PS2_CLK,
inout               PS2_DAT,

inout               PS2_CLK2,
inout               PS2_DAT2,

// Slider Switches
input       [ 9: 0] SW,

// Video-In
input               TD_CLK27,
input       [ 7: 0] TD_DATA,
input               TD_HS,
output              TD_RESET_N,
input               TD_VS,

// VGA
output      [ 7: 0] VGA_B,
output              VGA_BLANK_N,
output              VGA_CLK,
output      [ 7: 0] VGA_G,
output              VGA_HS,
output      [ 7: 0] VGA_R,
output              VGA_SYNC_N,
output              VGA_VS

);

//=======================================================
//  REG/WIRE declarations
//=======================================================

wire						system_clock;
wire						system_clock_locked;
wire						vga_clock;
wire						vga_clock_locked;

wire			[31: 0]	hex3_hex0;
wire			[15: 0]	hex5_hex4;

assign HEX0 = ~hex3_hex0[ 6: 0];
assign HEX1 = ~hex3_hex0[14: 8];
assign HEX2 = ~hex3_hex0[22:16];
assign HEX3 = ~hex3_hex0[30:24];
assign HEX4 = ~hex5_hex4[ 6: 0];
assign HEX5 = ~hex5_hex4[14: 8];

//=======================================================
//  Structural coding
//=======================================================

System_PLL_100 System_PLL (
	.refclk		(CLOCK_50),
	.rst			(1'b0),
	.outclk_0	(system_clock),
	.outclk_1	(DRAM_CLK),
	.locked		(system_clock_locked)
);

VGA_PLL VGA_PLL (
	.refclk		(CLOCK2_50),
	.rst			(1'b0),
	.outclk_0	(vga_clock),
	.locked		(vga_clock_locked)
);

Computer_System The_System (
	////////////////////////////////////
	// FPGA Side
	////////////////////////////////////

	// Global signals
	.sys_clk_ref_clk			(system_clock),
	.sys_clk_reset_n			(system_clock_locked),
	.vga_clk_ref_clk			(vga_clock),
	.vga_clk_reset_n			(1'b1),

    // ADC
	.adc_sclk							(ADC_SCLK),
	.adc_cs_n							(ADC_CONVST),
	.adc_dout							(ADC_SDO),
	.adc_din							(ADC_SDI),

	// AV Config
	.av_config_SCLK							(FPGA_I2C_SCLK),
	.av_config_SDAT							(FPGA_I2C_SDAT),

	// Audio Subsystem
	.audio_pll_ref_clk_clk					(CLOCK3_50),
	.audio_pll_ref_reset_reset				(1'b0),
	.audio_pll_clk_clk						(AUD_XCK),
	.audio_ADCDAT								(AUD_ADCDAT),
	.audio_ADCLRCK								(AUD_ADCLRCK),
	.audio_BCLK									(AUD_BCLK),
	.audio_DACDAT								(AUD_DACDAT),
	.audio_DACLRCK								(AUD_DACLRCK),

	// Slider Switches
	.slider_switches_export					(SW),

	// Pushbuttons
	.pushbuttons_export						(~KEY[3:0]),

	// Expansion JP1
    .expansion_jp1_export               ({GPIO[35:19], GPIO[17], GPIO[15:3], GPIO[1]}),

	// LEDs
	.leds_export								(LEDR),
	
	// Seven Segs
	.hex3_hex0_export							(hex3_hex0),
	.hex5_hex4_export							(hex5_hex4),
	
	// PS2 Ports
	.ps2_port_CLK								(PS2_CLK),
	.ps2_port_DAT								(PS2_DAT),
	.ps2_port_dual_CLK						(PS2_CLK2),
	.ps2_port_dual_DAT						(PS2_DAT2),

	// IrDA
	.irda_RXD									(IRDA_RXD),
	.irda_TXD									(IRDA_TXD),

	// VGA Subsystem
	.vga_CLK										(VGA_CLK),
	.vga_BLANK									(VGA_BLANK_N),
	.vga_SYNC									(VGA_SYNC_N),
	.vga_HS										(VGA_HS),
	.vga_VS										(VGA_VS),
	.vga_R										(VGA_R),
	.vga_G										(VGA_G),
	.vga_B										(VGA_B),
	
	// Video In Subsystem
	.video_in_TD_CLK27 						(TD_CLK27),
	.video_in_TD_DATA							(TD_DATA),
	.video_in_TD_HS							(TD_HS),
	.video_in_TD_VS							(TD_VS),
	.video_in_clk27_reset					(),
	.video_in_TD_RESET						(TD_RESET_N),
	.video_in_overflow_flag					(),
	
	// SDRAM
	.sdram_addr									(DRAM_ADDR),
	.sdram_ba									(DRAM_BA),
	.sdram_cas_n								(DRAM_CAS_N),
	.sdram_cke									(DRAM_CKE),
	.sdram_cs_n									(DRAM_CS_N),
	.sdram_dq									(DRAM_DQ),
	.sdram_dqm									({DRAM_UDQM,DRAM_LDQM}),
	.sdram_ras_n								(DRAM_RAS_N),
	.sdram_we_n									(DRAM_WE_N)
);


endmodule
